module sync_fifo_tb;
//testbench for sync fifo and alt sync fifo (Compare the results of sync fifo and alt sync fifo)

  endmodule