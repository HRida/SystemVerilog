// Class Definition
class MyFerrari;
  // Properties

  // Methods
  // Constructor
  function new(); //complete arguments
	  //complete here
  endfunction

  // Method to display information about the car
  function void displayInfo();
    $display(); //complete this 
  endfunction

  // Method to accelerate the car
  function void accelerate(); //add necessary argument
	  //complete here
  endfunction

  // Method to brake the car
  function void brake(); //add necessary argument
	  // complete here
  endfunction

endclass

