`ifndef DEFINES
`define DEFINES

`define NO_OF_TRANSACTIONS 100

`endif
 
