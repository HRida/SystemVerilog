`ifndef ADDER_4_BIT_DEFINES
`define ADDER_4_BIT_DEFINES


  `define ADDER_WIDTH 8
  `define NO_OF_TRANSACTIONS 1000

`endif
