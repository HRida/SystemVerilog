module dual_edge_detector (
  input logic clk,
  input logic reset,
  input logic signal,
  output logic pos_edge,
  output logic neg_edge
);

// .. your code goes here

endmodule
