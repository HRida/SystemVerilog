// Testbench
module MyFerrari_tb;
  // Instantiate the car object

  initial begin
    // Display initial information about the car
    // add code here
    
    // Accelerate the car
    // add code here

    // Brake the car
    // add code here

    // Display final information about the car
    // add code here

    // End simulation
    $finish;
  end
endmodule

